VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_bin_mult
  CLASS BLOCK ;
  FOREIGN wrapped_bin_mult ;
  ORIGIN 0.000 0.000 ;
  SIZE 220.000 BY 220.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 114.280 220.000 114.880 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 216.000 129.170 220.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 31.320 220.000 31.920 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 216.000 114.450 220.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 46.280 220.000 46.880 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 59.880 220.000 60.480 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 118.360 220.000 118.960 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 70.760 220.000 71.360 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 216.000 44.530 220.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 216.000 206.450 220.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 216.000 68.450 220.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 216.000 151.250 220.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 195.880 220.000 196.480 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 57.160 220.000 57.760 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 216.000 165.050 220.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 216.000 49.130 220.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 216.000 1.290 220.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 78.920 220.000 79.520 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 216.000 63.850 220.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 175.480 220.000 176.080 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 216.000 194.490 220.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 193.160 220.000 193.760 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 216.000 201.850 220.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 217.640 220.000 218.240 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 216.000 126.410 220.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.080 4.000 121.680 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 99.320 220.000 99.920 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 216.000 39.930 220.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 216.000 32.570 220.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 216.000 218.410 220.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 216.000 119.050 220.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 186.360 220.000 186.960 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 216.000 7.730 220.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 138.760 220.000 139.360 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 39.480 220.000 40.080 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 206.760 220.000 207.360 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 35.400 220.000 36.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 216.000 167.810 220.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 178.200 220.000 178.800 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 0.040 220.000 0.640 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 13.640 220.000 14.240 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.130 216.000 172.410 220.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 216.000 177.010 220.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 216.000 92.370 220.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 0.000 48.210 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 216.000 20.610 220.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 216.000 163.210 220.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 216.000 90.530 220.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 216.000 13.250 220.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 131.960 220.000 132.560 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 216.000 141.130 220.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 189.080 220.000 189.680 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 6.840 220.000 7.440 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 216.000 29.810 220.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 216.000 136.530 220.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 216.000 213.810 220.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 216.000 203.690 220.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 216.000 182.530 220.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 216.000 73.050 220.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 216.000 61.090 220.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 125.160 220.000 125.760 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 216.000 66.610 220.000 ;
    END
  END io_out[9]
  PIN rambus_wb_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END rambus_wb_ack_i
  PIN rambus_wb_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 156.440 220.000 157.040 ;
    END
  END rambus_wb_adr_o[0]
  PIN rambus_wb_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 216.000 15.090 220.000 ;
    END
  END rambus_wb_adr_o[1]
  PIN rambus_wb_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 216.000 75.810 220.000 ;
    END
  END rambus_wb_adr_o[2]
  PIN rambus_wb_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END rambus_wb_adr_o[3]
  PIN rambus_wb_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 214.920 220.000 215.520 ;
    END
  END rambus_wb_adr_o[4]
  PIN rambus_wb_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 42.200 220.000 42.800 ;
    END
  END rambus_wb_adr_o[5]
  PIN rambus_wb_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END rambus_wb_adr_o[6]
  PIN rambus_wb_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 103.400 220.000 104.000 ;
    END
  END rambus_wb_adr_o[7]
  PIN rambus_wb_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END rambus_wb_adr_o[8]
  PIN rambus_wb_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END rambus_wb_adr_o[9]
  PIN rambus_wb_clk_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END rambus_wb_clk_o
  PIN rambus_wb_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 216.000 53.730 220.000 ;
    END
  END rambus_wb_cyc_o
  PIN rambus_wb_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 216.000 85.930 220.000 ;
    END
  END rambus_wb_dat_i[0]
  PIN rambus_wb_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END rambus_wb_dat_i[10]
  PIN rambus_wb_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END rambus_wb_dat_i[11]
  PIN rambus_wb_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END rambus_wb_dat_i[12]
  PIN rambus_wb_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 21.800 220.000 22.400 ;
    END
  END rambus_wb_dat_i[13]
  PIN rambus_wb_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 216.000 117.210 220.000 ;
    END
  END rambus_wb_dat_i[14]
  PIN rambus_wb_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 216.000 83.170 220.000 ;
    END
  END rambus_wb_dat_i[15]
  PIN rambus_wb_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 216.000 102.490 220.000 ;
    END
  END rambus_wb_dat_i[16]
  PIN rambus_wb_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END rambus_wb_dat_i[17]
  PIN rambus_wb_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END rambus_wb_dat_i[18]
  PIN rambus_wb_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END rambus_wb_dat_i[19]
  PIN rambus_wb_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 0.000 31.650 4.000 ;
    END
  END rambus_wb_dat_i[1]
  PIN rambus_wb_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END rambus_wb_dat_i[20]
  PIN rambus_wb_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 216.000 95.130 220.000 ;
    END
  END rambus_wb_dat_i[21]
  PIN rambus_wb_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END rambus_wb_dat_i[22]
  PIN rambus_wb_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 110.200 220.000 110.800 ;
    END
  END rambus_wb_dat_i[23]
  PIN rambus_wb_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 121.080 220.000 121.680 ;
    END
  END rambus_wb_dat_i[24]
  PIN rambus_wb_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 149.640 220.000 150.240 ;
    END
  END rambus_wb_dat_i[25]
  PIN rambus_wb_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 216.000 124.570 220.000 ;
    END
  END rambus_wb_dat_i[26]
  PIN rambus_wb_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END rambus_wb_dat_i[27]
  PIN rambus_wb_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 216.000 34.410 220.000 ;
    END
  END rambus_wb_dat_i[28]
  PIN rambus_wb_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 167.320 220.000 167.920 ;
    END
  END rambus_wb_dat_i[29]
  PIN rambus_wb_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END rambus_wb_dat_i[2]
  PIN rambus_wb_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 2.760 220.000 3.360 ;
    END
  END rambus_wb_dat_i[30]
  PIN rambus_wb_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 216.000 87.770 220.000 ;
    END
  END rambus_wb_dat_i[31]
  PIN rambus_wb_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 107.480 220.000 108.080 ;
    END
  END rambus_wb_dat_i[3]
  PIN rambus_wb_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 74.840 220.000 75.440 ;
    END
  END rambus_wb_dat_i[4]
  PIN rambus_wb_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 216.000 17.850 220.000 ;
    END
  END rambus_wb_dat_i[5]
  PIN rambus_wb_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 216.000 51.890 220.000 ;
    END
  END rambus_wb_dat_i[6]
  PIN rambus_wb_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END rambus_wb_dat_i[7]
  PIN rambus_wb_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END rambus_wb_dat_i[8]
  PIN rambus_wb_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 216.000 184.370 220.000 ;
    END
  END rambus_wb_dat_i[9]
  PIN rambus_wb_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END rambus_wb_dat_o[0]
  PIN rambus_wb_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 4.000 ;
    END
  END rambus_wb_dat_o[10]
  PIN rambus_wb_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END rambus_wb_dat_o[11]
  PIN rambus_wb_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END rambus_wb_dat_o[12]
  PIN rambus_wb_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 127.880 220.000 128.480 ;
    END
  END rambus_wb_dat_o[13]
  PIN rambus_wb_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 216.000 27.050 220.000 ;
    END
  END rambus_wb_dat_o[14]
  PIN rambus_wb_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 216.000 191.730 220.000 ;
    END
  END rambus_wb_dat_o[15]
  PIN rambus_wb_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END rambus_wb_dat_o[16]
  PIN rambus_wb_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END rambus_wb_dat_o[17]
  PIN rambus_wb_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END rambus_wb_dat_o[18]
  PIN rambus_wb_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 216.000 111.690 220.000 ;
    END
  END rambus_wb_dat_o[19]
  PIN rambus_wb_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END rambus_wb_dat_o[1]
  PIN rambus_wb_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END rambus_wb_dat_o[20]
  PIN rambus_wb_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END rambus_wb_dat_o[21]
  PIN rambus_wb_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END rambus_wb_dat_o[22]
  PIN rambus_wb_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 53.080 220.000 53.680 ;
    END
  END rambus_wb_dat_o[23]
  PIN rambus_wb_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 216.000 148.490 220.000 ;
    END
  END rambus_wb_dat_o[24]
  PIN rambus_wb_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END rambus_wb_dat_o[25]
  PIN rambus_wb_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 216.000 121.810 220.000 ;
    END
  END rambus_wb_dat_o[26]
  PIN rambus_wb_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END rambus_wb_dat_o[27]
  PIN rambus_wb_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 210.840 220.000 211.440 ;
    END
  END rambus_wb_dat_o[28]
  PIN rambus_wb_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 216.000 22.450 220.000 ;
    END
  END rambus_wb_dat_o[29]
  PIN rambus_wb_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END rambus_wb_dat_o[2]
  PIN rambus_wb_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 164.600 220.000 165.200 ;
    END
  END rambus_wb_dat_o[30]
  PIN rambus_wb_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END rambus_wb_dat_o[31]
  PIN rambus_wb_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 216.000 99.730 220.000 ;
    END
  END rambus_wb_dat_o[3]
  PIN rambus_wb_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END rambus_wb_dat_o[4]
  PIN rambus_wb_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 216.000 153.090 220.000 ;
    END
  END rambus_wb_dat_o[5]
  PIN rambus_wb_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END rambus_wb_dat_o[6]
  PIN rambus_wb_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 24.520 220.000 25.120 ;
    END
  END rambus_wb_dat_o[7]
  PIN rambus_wb_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END rambus_wb_dat_o[8]
  PIN rambus_wb_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 216.000 80.410 220.000 ;
    END
  END rambus_wb_dat_o[9]
  PIN rambus_wb_rst_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END rambus_wb_rst_o
  PIN rambus_wb_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END rambus_wb_sel_o[0]
  PIN rambus_wb_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 216.000 155.850 220.000 ;
    END
  END rambus_wb_sel_o[1]
  PIN rambus_wb_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 216.000 71.210 220.000 ;
    END
  END rambus_wb_sel_o[2]
  PIN rambus_wb_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END rambus_wb_sel_o[3]
  PIN rambus_wb_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 216.000 145.730 220.000 ;
    END
  END rambus_wb_stb_o
  PIN rambus_wb_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END rambus_wb_we_o
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 206.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 206.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 206.960 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 216.000 133.770 220.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 216.000 175.170 220.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 216.000 109.850 220.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 216.000 59.250 220.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 96.600 220.000 97.200 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.610 216.000 5.890 220.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 216.000 199.090 220.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.160 4.000 125.760 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 216.000 107.090 220.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.610 216.000 143.890 220.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 68.040 220.000 68.640 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 160.520 220.000 161.120 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 216.000 216.570 220.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 28.600 220.000 29.200 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.770 216.000 211.050 220.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.210 216.000 10.490 220.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 216.000 131.930 220.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 146.920 220.000 147.520 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 216.000 37.170 220.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 216.000 46.370 220.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 216.000 41.770 220.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 63.960 220.000 64.560 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 216.000 189.890 220.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 204.040 220.000 204.640 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 216.000 78.570 220.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 85.720 220.000 86.320 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 199.960 220.000 200.560 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 136.040 220.000 136.640 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 216.000 209.210 220.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 216.000 105.250 220.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 92.520 220.000 93.120 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 10.920 220.000 11.520 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 50.360 220.000 50.960 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 216.000 197.250 220.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 171.400 220.000 172.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 89.800 220.000 90.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 182.280 220.000 182.880 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 216.000 187.130 220.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 0.000 200.930 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 216.000 179.770 220.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.720 4.000 154.320 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 216.000 138.370 220.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 216.000 97.890 220.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 216.000 170.570 220.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 17.720 220.000 18.320 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 153.720 220.000 154.320 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 142.840 220.000 143.440 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 216.000 160.450 220.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 216.000 157.690 220.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 216.000 25.210 220.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 216.000 56.490 220.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 216.000 3.130 220.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 216.000 81.640 220.000 82.240 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 7.225 217.895 215.135 ;
      LAYER met1 ;
        RECT 0.070 6.500 218.430 215.180 ;
      LAYER met2 ;
        RECT 0.100 215.720 0.730 218.125 ;
        RECT 1.570 215.720 2.570 218.125 ;
        RECT 3.410 215.720 5.330 218.125 ;
        RECT 6.170 215.720 7.170 218.125 ;
        RECT 8.010 215.720 9.930 218.125 ;
        RECT 10.770 215.720 12.690 218.125 ;
        RECT 13.530 215.720 14.530 218.125 ;
        RECT 15.370 215.720 17.290 218.125 ;
        RECT 18.130 215.720 20.050 218.125 ;
        RECT 20.890 215.720 21.890 218.125 ;
        RECT 22.730 215.720 24.650 218.125 ;
        RECT 25.490 215.720 26.490 218.125 ;
        RECT 27.330 215.720 29.250 218.125 ;
        RECT 30.090 215.720 32.010 218.125 ;
        RECT 32.850 215.720 33.850 218.125 ;
        RECT 34.690 215.720 36.610 218.125 ;
        RECT 37.450 215.720 39.370 218.125 ;
        RECT 40.210 215.720 41.210 218.125 ;
        RECT 42.050 215.720 43.970 218.125 ;
        RECT 44.810 215.720 45.810 218.125 ;
        RECT 46.650 215.720 48.570 218.125 ;
        RECT 49.410 215.720 51.330 218.125 ;
        RECT 52.170 215.720 53.170 218.125 ;
        RECT 54.010 215.720 55.930 218.125 ;
        RECT 56.770 215.720 58.690 218.125 ;
        RECT 59.530 215.720 60.530 218.125 ;
        RECT 61.370 215.720 63.290 218.125 ;
        RECT 64.130 215.720 66.050 218.125 ;
        RECT 66.890 215.720 67.890 218.125 ;
        RECT 68.730 215.720 70.650 218.125 ;
        RECT 71.490 215.720 72.490 218.125 ;
        RECT 73.330 215.720 75.250 218.125 ;
        RECT 76.090 215.720 78.010 218.125 ;
        RECT 78.850 215.720 79.850 218.125 ;
        RECT 80.690 215.720 82.610 218.125 ;
        RECT 83.450 215.720 85.370 218.125 ;
        RECT 86.210 215.720 87.210 218.125 ;
        RECT 88.050 215.720 89.970 218.125 ;
        RECT 90.810 215.720 91.810 218.125 ;
        RECT 92.650 215.720 94.570 218.125 ;
        RECT 95.410 215.720 97.330 218.125 ;
        RECT 98.170 215.720 99.170 218.125 ;
        RECT 100.010 215.720 101.930 218.125 ;
        RECT 102.770 215.720 104.690 218.125 ;
        RECT 105.530 215.720 106.530 218.125 ;
        RECT 107.370 215.720 109.290 218.125 ;
        RECT 110.130 215.720 111.130 218.125 ;
        RECT 111.970 215.720 113.890 218.125 ;
        RECT 114.730 215.720 116.650 218.125 ;
        RECT 117.490 215.720 118.490 218.125 ;
        RECT 119.330 215.720 121.250 218.125 ;
        RECT 122.090 215.720 124.010 218.125 ;
        RECT 124.850 215.720 125.850 218.125 ;
        RECT 126.690 215.720 128.610 218.125 ;
        RECT 129.450 215.720 131.370 218.125 ;
        RECT 132.210 215.720 133.210 218.125 ;
        RECT 134.050 215.720 135.970 218.125 ;
        RECT 136.810 215.720 137.810 218.125 ;
        RECT 138.650 215.720 140.570 218.125 ;
        RECT 141.410 215.720 143.330 218.125 ;
        RECT 144.170 215.720 145.170 218.125 ;
        RECT 146.010 215.720 147.930 218.125 ;
        RECT 148.770 215.720 150.690 218.125 ;
        RECT 151.530 215.720 152.530 218.125 ;
        RECT 153.370 215.720 155.290 218.125 ;
        RECT 156.130 215.720 157.130 218.125 ;
        RECT 157.970 215.720 159.890 218.125 ;
        RECT 160.730 215.720 162.650 218.125 ;
        RECT 163.490 215.720 164.490 218.125 ;
        RECT 165.330 215.720 167.250 218.125 ;
        RECT 168.090 215.720 170.010 218.125 ;
        RECT 170.850 215.720 171.850 218.125 ;
        RECT 172.690 215.720 174.610 218.125 ;
        RECT 175.450 215.720 176.450 218.125 ;
        RECT 177.290 215.720 179.210 218.125 ;
        RECT 180.050 215.720 181.970 218.125 ;
        RECT 182.810 215.720 183.810 218.125 ;
        RECT 184.650 215.720 186.570 218.125 ;
        RECT 187.410 215.720 189.330 218.125 ;
        RECT 190.170 215.720 191.170 218.125 ;
        RECT 192.010 215.720 193.930 218.125 ;
        RECT 194.770 215.720 196.690 218.125 ;
        RECT 197.530 215.720 198.530 218.125 ;
        RECT 199.370 215.720 201.290 218.125 ;
        RECT 202.130 215.720 203.130 218.125 ;
        RECT 203.970 215.720 205.890 218.125 ;
        RECT 206.730 215.720 208.650 218.125 ;
        RECT 209.490 215.720 210.490 218.125 ;
        RECT 211.330 215.720 213.250 218.125 ;
        RECT 214.090 215.720 216.010 218.125 ;
        RECT 216.850 215.720 217.850 218.125 ;
        RECT 0.100 4.280 218.400 215.720 ;
        RECT 0.650 0.155 1.650 4.280 ;
        RECT 2.490 0.155 4.410 4.280 ;
        RECT 5.250 0.155 6.250 4.280 ;
        RECT 7.090 0.155 9.010 4.280 ;
        RECT 9.850 0.155 11.770 4.280 ;
        RECT 12.610 0.155 13.610 4.280 ;
        RECT 14.450 0.155 16.370 4.280 ;
        RECT 17.210 0.155 19.130 4.280 ;
        RECT 19.970 0.155 20.970 4.280 ;
        RECT 21.810 0.155 23.730 4.280 ;
        RECT 24.570 0.155 25.570 4.280 ;
        RECT 26.410 0.155 28.330 4.280 ;
        RECT 29.170 0.155 31.090 4.280 ;
        RECT 31.930 0.155 32.930 4.280 ;
        RECT 33.770 0.155 35.690 4.280 ;
        RECT 36.530 0.155 38.450 4.280 ;
        RECT 39.290 0.155 40.290 4.280 ;
        RECT 41.130 0.155 43.050 4.280 ;
        RECT 43.890 0.155 44.890 4.280 ;
        RECT 45.730 0.155 47.650 4.280 ;
        RECT 48.490 0.155 50.410 4.280 ;
        RECT 51.250 0.155 52.250 4.280 ;
        RECT 53.090 0.155 55.010 4.280 ;
        RECT 55.850 0.155 57.770 4.280 ;
        RECT 58.610 0.155 59.610 4.280 ;
        RECT 60.450 0.155 62.370 4.280 ;
        RECT 63.210 0.155 64.210 4.280 ;
        RECT 65.050 0.155 66.970 4.280 ;
        RECT 67.810 0.155 69.730 4.280 ;
        RECT 70.570 0.155 71.570 4.280 ;
        RECT 72.410 0.155 74.330 4.280 ;
        RECT 75.170 0.155 77.090 4.280 ;
        RECT 77.930 0.155 78.930 4.280 ;
        RECT 79.770 0.155 81.690 4.280 ;
        RECT 82.530 0.155 84.450 4.280 ;
        RECT 85.290 0.155 86.290 4.280 ;
        RECT 87.130 0.155 89.050 4.280 ;
        RECT 89.890 0.155 90.890 4.280 ;
        RECT 91.730 0.155 93.650 4.280 ;
        RECT 94.490 0.155 96.410 4.280 ;
        RECT 97.250 0.155 98.250 4.280 ;
        RECT 99.090 0.155 101.010 4.280 ;
        RECT 101.850 0.155 103.770 4.280 ;
        RECT 104.610 0.155 105.610 4.280 ;
        RECT 106.450 0.155 108.370 4.280 ;
        RECT 109.210 0.155 110.210 4.280 ;
        RECT 111.050 0.155 112.970 4.280 ;
        RECT 113.810 0.155 115.730 4.280 ;
        RECT 116.570 0.155 117.570 4.280 ;
        RECT 118.410 0.155 120.330 4.280 ;
        RECT 121.170 0.155 123.090 4.280 ;
        RECT 123.930 0.155 124.930 4.280 ;
        RECT 125.770 0.155 127.690 4.280 ;
        RECT 128.530 0.155 129.530 4.280 ;
        RECT 130.370 0.155 132.290 4.280 ;
        RECT 133.130 0.155 135.050 4.280 ;
        RECT 135.890 0.155 136.890 4.280 ;
        RECT 137.730 0.155 139.650 4.280 ;
        RECT 140.490 0.155 142.410 4.280 ;
        RECT 143.250 0.155 144.250 4.280 ;
        RECT 145.090 0.155 147.010 4.280 ;
        RECT 147.850 0.155 149.770 4.280 ;
        RECT 150.610 0.155 151.610 4.280 ;
        RECT 152.450 0.155 154.370 4.280 ;
        RECT 155.210 0.155 156.210 4.280 ;
        RECT 157.050 0.155 158.970 4.280 ;
        RECT 159.810 0.155 161.730 4.280 ;
        RECT 162.570 0.155 163.570 4.280 ;
        RECT 164.410 0.155 166.330 4.280 ;
        RECT 167.170 0.155 169.090 4.280 ;
        RECT 169.930 0.155 170.930 4.280 ;
        RECT 171.770 0.155 173.690 4.280 ;
        RECT 174.530 0.155 175.530 4.280 ;
        RECT 176.370 0.155 178.290 4.280 ;
        RECT 179.130 0.155 181.050 4.280 ;
        RECT 181.890 0.155 182.890 4.280 ;
        RECT 183.730 0.155 185.650 4.280 ;
        RECT 186.490 0.155 188.410 4.280 ;
        RECT 189.250 0.155 190.250 4.280 ;
        RECT 191.090 0.155 193.010 4.280 ;
        RECT 193.850 0.155 194.850 4.280 ;
        RECT 195.690 0.155 197.610 4.280 ;
        RECT 198.450 0.155 200.370 4.280 ;
        RECT 201.210 0.155 202.210 4.280 ;
        RECT 203.050 0.155 204.970 4.280 ;
        RECT 205.810 0.155 207.730 4.280 ;
        RECT 208.570 0.155 209.570 4.280 ;
        RECT 210.410 0.155 212.330 4.280 ;
        RECT 213.170 0.155 215.090 4.280 ;
        RECT 215.930 0.155 216.930 4.280 ;
        RECT 217.770 0.155 218.400 4.280 ;
      LAYER met3 ;
        RECT 4.400 217.240 215.600 218.105 ;
        RECT 4.000 215.920 216.000 217.240 ;
        RECT 4.000 214.560 215.600 215.920 ;
        RECT 4.400 214.520 215.600 214.560 ;
        RECT 4.400 213.160 216.000 214.520 ;
        RECT 4.000 211.840 216.000 213.160 ;
        RECT 4.400 210.440 215.600 211.840 ;
        RECT 4.000 207.760 216.000 210.440 ;
        RECT 4.400 206.360 215.600 207.760 ;
        RECT 4.000 205.040 216.000 206.360 ;
        RECT 4.000 203.680 215.600 205.040 ;
        RECT 4.400 203.640 215.600 203.680 ;
        RECT 4.400 202.280 216.000 203.640 ;
        RECT 4.000 200.960 216.000 202.280 ;
        RECT 4.400 199.560 215.600 200.960 ;
        RECT 4.000 196.880 216.000 199.560 ;
        RECT 4.400 195.480 215.600 196.880 ;
        RECT 4.000 194.160 216.000 195.480 ;
        RECT 4.000 192.800 215.600 194.160 ;
        RECT 4.400 192.760 215.600 192.800 ;
        RECT 4.400 191.400 216.000 192.760 ;
        RECT 4.000 190.080 216.000 191.400 ;
        RECT 4.400 188.680 215.600 190.080 ;
        RECT 4.000 187.360 216.000 188.680 ;
        RECT 4.000 186.000 215.600 187.360 ;
        RECT 4.400 185.960 215.600 186.000 ;
        RECT 4.400 184.600 216.000 185.960 ;
        RECT 4.000 183.280 216.000 184.600 ;
        RECT 4.400 181.880 215.600 183.280 ;
        RECT 4.000 179.200 216.000 181.880 ;
        RECT 4.400 177.800 215.600 179.200 ;
        RECT 4.000 176.480 216.000 177.800 ;
        RECT 4.000 175.120 215.600 176.480 ;
        RECT 4.400 175.080 215.600 175.120 ;
        RECT 4.400 173.720 216.000 175.080 ;
        RECT 4.000 172.400 216.000 173.720 ;
        RECT 4.400 171.000 215.600 172.400 ;
        RECT 4.000 168.320 216.000 171.000 ;
        RECT 4.400 166.920 215.600 168.320 ;
        RECT 4.000 165.600 216.000 166.920 ;
        RECT 4.000 164.240 215.600 165.600 ;
        RECT 4.400 164.200 215.600 164.240 ;
        RECT 4.400 162.840 216.000 164.200 ;
        RECT 4.000 161.520 216.000 162.840 ;
        RECT 4.400 160.120 215.600 161.520 ;
        RECT 4.000 157.440 216.000 160.120 ;
        RECT 4.400 156.040 215.600 157.440 ;
        RECT 4.000 154.720 216.000 156.040 ;
        RECT 4.400 153.320 215.600 154.720 ;
        RECT 4.000 150.640 216.000 153.320 ;
        RECT 4.400 149.240 215.600 150.640 ;
        RECT 4.000 147.920 216.000 149.240 ;
        RECT 4.000 146.560 215.600 147.920 ;
        RECT 4.400 146.520 215.600 146.560 ;
        RECT 4.400 145.160 216.000 146.520 ;
        RECT 4.000 143.840 216.000 145.160 ;
        RECT 4.400 142.440 215.600 143.840 ;
        RECT 4.000 139.760 216.000 142.440 ;
        RECT 4.400 138.360 215.600 139.760 ;
        RECT 4.000 137.040 216.000 138.360 ;
        RECT 4.000 135.680 215.600 137.040 ;
        RECT 4.400 135.640 215.600 135.680 ;
        RECT 4.400 134.280 216.000 135.640 ;
        RECT 4.000 132.960 216.000 134.280 ;
        RECT 4.400 131.560 215.600 132.960 ;
        RECT 4.000 128.880 216.000 131.560 ;
        RECT 4.400 127.480 215.600 128.880 ;
        RECT 4.000 126.160 216.000 127.480 ;
        RECT 4.400 124.760 215.600 126.160 ;
        RECT 4.000 122.080 216.000 124.760 ;
        RECT 4.400 120.680 215.600 122.080 ;
        RECT 4.000 119.360 216.000 120.680 ;
        RECT 4.000 118.000 215.600 119.360 ;
        RECT 4.400 117.960 215.600 118.000 ;
        RECT 4.400 116.600 216.000 117.960 ;
        RECT 4.000 115.280 216.000 116.600 ;
        RECT 4.400 113.880 215.600 115.280 ;
        RECT 4.000 111.200 216.000 113.880 ;
        RECT 4.400 109.800 215.600 111.200 ;
        RECT 4.000 108.480 216.000 109.800 ;
        RECT 4.000 107.120 215.600 108.480 ;
        RECT 4.400 107.080 215.600 107.120 ;
        RECT 4.400 105.720 216.000 107.080 ;
        RECT 4.000 104.400 216.000 105.720 ;
        RECT 4.400 103.000 215.600 104.400 ;
        RECT 4.000 100.320 216.000 103.000 ;
        RECT 4.400 98.920 215.600 100.320 ;
        RECT 4.000 97.600 216.000 98.920 ;
        RECT 4.000 96.240 215.600 97.600 ;
        RECT 4.400 96.200 215.600 96.240 ;
        RECT 4.400 94.840 216.000 96.200 ;
        RECT 4.000 93.520 216.000 94.840 ;
        RECT 4.400 92.120 215.600 93.520 ;
        RECT 4.000 90.800 216.000 92.120 ;
        RECT 4.000 89.440 215.600 90.800 ;
        RECT 4.400 89.400 215.600 89.440 ;
        RECT 4.400 88.040 216.000 89.400 ;
        RECT 4.000 86.720 216.000 88.040 ;
        RECT 4.400 85.320 215.600 86.720 ;
        RECT 4.000 82.640 216.000 85.320 ;
        RECT 4.400 81.240 215.600 82.640 ;
        RECT 4.000 79.920 216.000 81.240 ;
        RECT 4.000 78.560 215.600 79.920 ;
        RECT 4.400 78.520 215.600 78.560 ;
        RECT 4.400 77.160 216.000 78.520 ;
        RECT 4.000 75.840 216.000 77.160 ;
        RECT 4.400 74.440 215.600 75.840 ;
        RECT 4.000 71.760 216.000 74.440 ;
        RECT 4.400 70.360 215.600 71.760 ;
        RECT 4.000 69.040 216.000 70.360 ;
        RECT 4.000 67.680 215.600 69.040 ;
        RECT 4.400 67.640 215.600 67.680 ;
        RECT 4.400 66.280 216.000 67.640 ;
        RECT 4.000 64.960 216.000 66.280 ;
        RECT 4.400 63.560 215.600 64.960 ;
        RECT 4.000 60.880 216.000 63.560 ;
        RECT 4.400 59.480 215.600 60.880 ;
        RECT 4.000 58.160 216.000 59.480 ;
        RECT 4.400 56.760 215.600 58.160 ;
        RECT 4.000 54.080 216.000 56.760 ;
        RECT 4.400 52.680 215.600 54.080 ;
        RECT 4.000 51.360 216.000 52.680 ;
        RECT 4.000 50.000 215.600 51.360 ;
        RECT 4.400 49.960 215.600 50.000 ;
        RECT 4.400 48.600 216.000 49.960 ;
        RECT 4.000 47.280 216.000 48.600 ;
        RECT 4.400 45.880 215.600 47.280 ;
        RECT 4.000 43.200 216.000 45.880 ;
        RECT 4.400 41.800 215.600 43.200 ;
        RECT 4.000 40.480 216.000 41.800 ;
        RECT 4.000 39.120 215.600 40.480 ;
        RECT 4.400 39.080 215.600 39.120 ;
        RECT 4.400 37.720 216.000 39.080 ;
        RECT 4.000 36.400 216.000 37.720 ;
        RECT 4.400 35.000 215.600 36.400 ;
        RECT 4.000 32.320 216.000 35.000 ;
        RECT 4.400 30.920 215.600 32.320 ;
        RECT 4.000 29.600 216.000 30.920 ;
        RECT 4.400 28.200 215.600 29.600 ;
        RECT 4.000 25.520 216.000 28.200 ;
        RECT 4.400 24.120 215.600 25.520 ;
        RECT 4.000 22.800 216.000 24.120 ;
        RECT 4.000 21.440 215.600 22.800 ;
        RECT 4.400 21.400 215.600 21.440 ;
        RECT 4.400 20.040 216.000 21.400 ;
        RECT 4.000 18.720 216.000 20.040 ;
        RECT 4.400 17.320 215.600 18.720 ;
        RECT 4.000 14.640 216.000 17.320 ;
        RECT 4.400 13.240 215.600 14.640 ;
        RECT 4.000 11.920 216.000 13.240 ;
        RECT 4.000 10.560 215.600 11.920 ;
        RECT 4.400 10.520 215.600 10.560 ;
        RECT 4.400 9.160 216.000 10.520 ;
        RECT 4.000 7.840 216.000 9.160 ;
        RECT 4.400 6.440 215.600 7.840 ;
        RECT 4.000 3.760 216.000 6.440 ;
        RECT 4.400 2.360 215.600 3.760 ;
        RECT 4.000 1.040 216.000 2.360 ;
        RECT 4.000 0.175 215.600 1.040 ;
      LAYER met4 ;
        RECT 116.215 80.415 116.545 92.985 ;
  END
END wrapped_bin_mult
END LIBRARY

